Template: debian-installer/main-menu
Type: select
Choices: ${MENU}
Choices-sv: ${MENU}
Default: ${DEFAULT}
Description: Choose the next step:
 Here is the main menu of the Debian installer.
Description-sv: Välj nästa steg:
 Det här är huvudmenyn för Debians installationsprogram.
