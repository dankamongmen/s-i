Template: anna/retriever
Type: select
Choices: ${CHOICES}
Choices-sv: ${CHOICES}
Default: ${DEFAULT}
Default-sv: ${DEFAULT}
Description: Choose the retriever to use.
 The retriever is responsible for fetching the packages to be
 installed.
Description-sv: V�lj vilken h�mtare (retriever) som ska anv�ndas.
 H�mtaren ansvarar f�r att h�mta paketen som ska installeras.
